library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Li_Memory is

	port(
		clk: in std_logic;
		read_address: in std_logic_vector(31 downto 0);
		data: in std_logic_vector(31 downto 0);
		wren, rd: in std_logic;
		q: out std_logic_vector(31 downto 0)
	);
	
end Li_Memory;

architecture arch of Li_Memory is

	signal ram_addr: std_logic_vector(31 downto 0);
	type data_memory is array (0 to 31) of std_logic_vector(31 downto 0);
	signal ram: data_memory := (
		"00000000000000000000000000001010", -- 10
		"00000000000000000000000000010100", -- 20
		"00000000000000000000000000011110", -- 30
		"00000000000000000000000000101000", -- 40
		"00000000000000000000000000110010", -- 50
		"00000000000000000000000000111100", -- 60
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000",
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000", 
		"00000000000000000000000000000000"
		
	);
	
	begin
	
		ram_addr <= ram_addr(31 downto 0);
		process(clk)
			begin
				if(rising_edge(clk)) then
					if(wren = '1') then
					ram(to_integer(unsigned(ram_addr))) <= data;
					end if;
				end if;
		end process;
				
		q <= ram(to_integer(unsigned(ram_addr))) when (rd = '1') else x"00000000";
		
end arch;
					
					
					
					
		